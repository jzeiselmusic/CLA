module final_test_bench();

	logic [15:0] A0;
	logic [15:0] B0;
	logic [15:0] SUM0;
	logic [15:0] DIFF0;
	logic [15:0] ABS0;
	logic S_OF0;
	logic D_OF0;
	logic LT0;

	top_level ALU(A0[15:0], B0[15:0], SUM0[15:0], 
		DIFF0[15:0], ABS0[15:0], S_OF0, D_OF0, LT0);

	initial begin

		A0 = 16'b0110110000111100;  
		B0 = 16'b0000000000110000; 
		#100;

		//SUM should be 0110110001101100 // 27756
		//ABS should be 0110110001101100 // 27756

		A0 = 16'b1111111100111000;
		B0 = 16'b1111110000011000;
		#100;

		//SUM should be 1111101101010000 // -1200
		//ABS should be 0000010010110000 // 1200

		A0 = 16'b0001001110001000;
		B0 = 16'b0111100100011000;
		#100;
		
		// SUM IS INCORRECT
		// S_OF is 1

		A0 = 16'b1000011011101000;
		B0 = 16'b1110110001111000;
		#100;
		
		// SUM IS INCORRECT 
		// S_OF is 1

		A0 = 16'b0111100100011000;
		B0 = 16'b1110110001111000;
		#100;

		// SUM should be 0110010110010000 // 26000
		// ABS should be 0110010110010000 // 26000

		A0 = 16'b1111111100111000;
		B0 = 16'b0000000111110100;
		#100;

		//SUM should be 0000000100101100 // 300
		//ABS should be 0000000100101100 // 300

		A0 = 16'b0000000011001000;
		B0 = 16'b1111111000001100;
		#100;

		// SUM should be 1111111011010100 // -300
		// ABS should be 0000000100101100 // 300

		A0 = 16'b1000011011101000;
		B0 = 16'b0001001110001000;

		//SUM should be 1001101001110000 // -26000
		//ABS should be 0110010110010000 // 26000

	end

endmodule
